`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: An-Ting Hsu
// 
// Create Date:    03:45:20 05/22/2015 
// Module Name:    music 
// Project Name:   Lab10-2
// Revision: 
// Revision 0.01 - File Created
//
//////////////////////////////////////////////////////////////////////////////////
`define BIT_WIDTH 10
module music(
	q0, //shifter output
	clk, // global clock
	rst_n //active low reset
);

output reg [`BIT_WIDTH-1:0] q0; //output
reg [`BIT_WIDTH-1:0] q1, q2, q3, q4, q5, q6, q7, q8, q9;
reg [`BIT_WIDTH-1:0] q10, q11, q12, q13, q14, q15, q16, q17, q18, q19;
reg [`BIT_WIDTH-1:0] q20, q21, q22, q23, q24, q25, q26, q27, q28, q29;
reg [`BIT_WIDTH-1:0] q30, q31, q32, q33, q34, q35, q36, q37, q38, q39;
reg [`BIT_WIDTH-1:0] q40, q41, q42, q43, q44, q45, q46, q47, q48, q49;
reg [`BIT_WIDTH-1:0] q50, q51, q52, q53, q54, q55, q56, q57, q58, q59;
reg [`BIT_WIDTH-1:0] q60, q61, q62, q63, q64, q65, q66, q67, q68, q69;
reg [`BIT_WIDTH-1:0] q70, q71, q72, q73, q74, q75, q76, q77, q78, q79;
reg [`BIT_WIDTH-1:0] q80, q81, q82, q83, q84, q85, q86, q87, q88, q89;
reg [`BIT_WIDTH-1:0] q90, q91, q92, q93, q94, q95, q96, q97, q98, q99;
reg [`BIT_WIDTH-1:0] q100, q101, q102, q103, q104, q105, q106, q107, q108, q109;
reg [`BIT_WIDTH-1:0] q110, q111, q112, q113, q114, q115, q116, q117, q118, q119;
reg [`BIT_WIDTH-1:0] q120, q121, q122, q123, q124, q125, q126, q127, q128, q129;
reg [`BIT_WIDTH-1:0] q130, q131, q132;
input clk, rst_n; //clock & global clock

//Sequential logics: Flip Flops
always @(posedge clk or negedge rst_n)
	if(~rst_n)
		begin
			q0 <= {6'd47, 4'd0};
			q1 <= {6'd15, 4'd2};
			q2 <= {6'd15, 4'd5};
			q3 <= {6'd7, 4'd4};
			q4 <= {6'd7, 4'd5};
			q5 <= {6'd15, 4'd6};
			q6 <= {6'd7, 4'd5};
			q7 <= {6'd7, 4'd6};
			q8 <= {6'd7, 4'd7};
			q9 <= {6'd7, 4'd7};
			q10 <= {6'd7, 4'd8};
			q11 <= {6'd7, 4'd7};
			q12 <= {6'd15, 4'd3};
			q13 <= {6'd7, 4'd6};
			q14 <= {6'd7, 4'd6};
			q15 <= {6'd15, 4'd5};
			q16 <= {6'd7, 4'd5};
			q17 <= {6'd7, 4'd5};
			q18 <= {6'd15, 4'd4};
			q19 <= {6'd7, 4'd3};
			q20 <= {6'd7, 4'd4};
			q21 <= {6'd47, 4'd5};
			q22 <= {6'd15, 4'd2};
			q23 <= {6'd15, 4'd5};
			q24 <= {6'd7, 4'd4};
			q25 <= {6'd7, 4'd5};
			q26 <= {6'd15, 4'd6};
			q27 <= {6'd7, 4'd5};
			q28 <= {6'd7, 4'd6};
			q29 <= {6'd7, 4'd7};
			q30 <= {6'd7, 4'd7};
			q31 <= {6'd7, 4'd8};
			q32 <= {6'd7, 4'd7};
			q33 <= {6'd15, 4'd3};
			q34 <= {6'd7, 4'd6};
			q35 <= {6'd7, 4'd6};
			q36 <= {6'd15, 4'd5};
			q37 <= {6'd7, 4'd5};
			q38 <= {6'd7, 4'd5};
			q39 <= {6'd15, 4'd4};
			q40 <= {6'd7, 4'd3};
			q41 <= {6'd7, 4'd4};
			q42 <= {6'd47, 4'd5};
			q43 <= {6'd7, 4'd5};
			q44 <= {6'd7, 4'd7};
			q45 <= {6'd15, 4'd9};
			q46 <= {6'd7, 4'd7};
			q47 <= {6'd7, 4'd6};
			q48 <= {6'd15, 4'd5};
			q49 <= {6'd7, 4'd4};
			q50 <= {6'd7, 4'd5};
			q51 <= {6'd7, 4'd6};
			q52 <= {6'd7, 4'd5};
			q53 <= {6'd7, 4'd4};
			q54 <= {6'd7, 4'd3};
			q55 <= {6'd15, 4'd2};
			q56 <= {6'd7, 4'd5};
			q57 <= {6'd7, 4'd7};
			q58 <= {6'd15, 4'd9};
			q59 <= {6'd7, 4'd7};
			q60 <= {6'd7, 4'd6};
			q61 <= {6'd7, 4'd5};
			q62 <= {6'd3, 4'd6};
			q63 <= {6'd3, 4'd5};
			q64 <= {6'd7, 4'd4};
			q65 <= {6'd7, 4'd5};
			q66 <= {6'd47, 4'd6};
			q67 <= {6'd7, 4'd0};
			q68 <= {6'd7, 4'd2};
			q69 <= {6'd7, 4'd5};
			q70 <= {6'd7, 4'd5};
			q71 <= {6'd15, 4'd0};
			q72 <= {6'd7, 4'd6};
			q73 <= {6'd15, 4'd6};
			q74 <= {6'd7, 4'd0};
			q75 <= {6'd7, 4'd7};
			q76 <= {6'd7, 4'd7};
			q77 <= {6'd7, 4'd8};
			q78 <= {6'd7, 4'd7};
			q79 <= {6'd15, 4'd3};
			q80 <= {6'd7, 4'd6};
			q81 <= {6'd7, 4'd6};
			q82 <= {6'd15, 4'd5};
			q83 <= {6'd7, 4'd5};
			q84 <= {6'd7, 4'd5};
			q85 <= {6'd15, 4'd4};
			q86 <= {6'd7, 4'd3};
			q87 <= {6'd7, 4'd4};
			q88 <= {6'd47, 4'd5};
			q89 <= {6'd15, 4'd2};
			q90 <= {6'd15, 4'd5};
			q91 <= {6'd7, 4'd2};
			q92 <= {6'd7, 4'd2};
			q93 <= {6'd7, 4'd3};
			q94 <= {6'd7, 4'd3};
			q95 <= {6'd15, 4'd2};
			q96 <= {6'd15, 4'd1};
			q97 <= {6'd15, 4'd2};
			q98 <= {6'd15, 4'd1};
			q99 <= {6'd7, 4'd2};
			q100 <= {6'd7, 4'd2};
			q101 <= {6'd15, 4'd5};
			q102 <= {6'd7, 4'd2};
			q103 <= {6'd7, 4'd2};
			q104 <= {6'd7, 4'd3};
			q105 <= {6'd7, 4'd3};
			q106 <= {6'd15, 4'd2};
			q107 <= {6'd15, 4'd1};
			q108 <= {6'd15, 4'd2};
			q109 <= {6'd15, 4'd1};
			q110 <= {6'd7, 4'd2};
			q111 <= {6'd7, 4'd2};
			q112 <= {6'd7, 4'd5};
			q113 <= {6'd7, 4'd5};
			q114 <= {6'd15, 4'd0};
			q115 <= {6'd7, 4'd6};
			q116 <= {6'd15, 4'd6};
			q117 <= {6'd7, 4'd0};
			q118 <= {6'd7, 4'd7};
			q119 <= {6'd7, 4'd7};
			q120 <= {6'd7, 4'd8};
			q121 <= {6'd7, 4'd7};
			q122 <= {6'd15, 4'd3};
			q123 <= {6'd7, 4'd6};
			q124 <= {6'd7, 4'd6};
			q125 <= {6'd15, 4'd5};
			q126 <= {6'd15, 4'd4};
			q127 <= {6'd7, 4'd3};
			q128 <= {6'd7, 4'd4};
			q129 <= {6'd15, 4'd5};
			q130 <= {6'd15, 4'd0};
			q131 <= {6'd71, 4'd0};
			q132 <= {6'd71, 4'd0};
		end
	else
		begin
			q0 <= q1;
			q1 <= q2;
			q2 <= q3;
			q3 <= q4;
			q4 <= q5;
			q5 <= q6;
			q6 <= q7;
			q7 <= q8;
			q8 <= q9;
			q9 <= q10;
			q10 <= q11;
			q11 <= q12;
			q12 <= q13;
			q13 <= q14;
			q14 <= q15;
			q15 <= q16;
			q16 <= q17;
			q17 <= q18;
			q18 <= q19;
			q19 <= q20;
			q20 <= q21;
			q21 <= q22;
			q22 <= q23;
			q23 <= q24;
			q24 <= q25;
			q25 <= q26;
			q26 <= q27;
			q27 <= q28;
			q28 <= q29;
			q29 <= q30;
			q30 <= q31;
			q31 <= q32;
			q32 <= q33;
			q33 <= q34;
			q34 <= q35;
			q35 <= q36;
			q36 <= q37;
			q37 <= q38;
			q38 <= q39;
			q39 <= q40;
			q40 <= q41;
			q41 <= q42;
			q42 <= q43;
			q43 <= q44;
			q44 <= q45;
			q45 <= q46;
			q46 <= q47;
			q47 <= q48;
			q48 <= q49;
			q49 <= q50;
			q50 <= q51;
			q51 <= q52;
			q52 <= q53;
			q53 <= q54;
			q54 <= q55;
			q55 <= q56;
			q56 <= q57;
			q57 <= q58;
			q58 <= q59;
			q59 <= q60;
			q60 <= q61;
			q61 <= q62;
			q62 <= q63;
			q63 <= q64;
			q64 <= q65;
			q65 <= q66;
			q66 <= q67;
			q67 <= q68;
			q68 <= q69;
			q69 <= q70;
			q70 <= q71;
			q71 <= q72;
			q72 <= q73;
			q73 <= q74;
			q74 <= q75;
			q75 <= q76;
			q76 <= q77;
			q77 <= q78;
			q78 <= q79;
			q79 <= q80;
			q80 <= q81;
			q81 <= q82;
			q82 <= q83;
			q83 <= q84;
			q84 <= q85;
			q85 <= q86;
			q86 <= q87;
			q87 <= q88;
			q88 <= q89;
			q89 <= q90;
			q90 <= q91;
			q91 <= q92;
			q92 <= q93;
			q93 <= q94;
			q94 <= q95;
			q95 <= q96;
			q96 <= q97;
			q97 <= q98;
			q98 <= q99;
			q99 <= q100;
			q100 <= q101;
			q101 <= q102;
			q102 <= q103;
			q103 <= q104;
			q104 <= q105;
			q105 <= q106;
			q106 <= q107;
			q107 <= q108;
			q108 <= q109;
			q109 <= q110;
			q110 <= q111;
			q111 <= q112;
			q112 <= q113;
			q113 <= q114;
			q114 <= q115;
			q115 <= q116;
			q116 <= q117;
			q117 <= q118;
			q118 <= q119;
			q119 <= q120;
			q120 <= q121;
			q121 <= q122;
			q122 <= q123;
			q123 <= q124;
			q124 <= q125;
			q125 <= q126;
			q126 <= q127;
			q127 <= q128;
			q128 <= q129;
			q129 <= q130;
			q130 <= q131;
			q131 <= q132;
			q132 <= q0;
		end
endmodule
